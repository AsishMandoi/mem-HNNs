*HNN_proj

.MODEL NMOS

M1SSL BL1 G01 S11 S11 NMOS
M11 S11 G11 S21 S21 NMOS
M21 S21 G21 S31 S31 NMOS
M31 S31 G31 S41 S41 NMOS
M41 S41 G41 S51 S51 NMOS

M2SSL BL2 G02 S12 S12 NMOS
M12 S12 G12 S22 S22 NMOS
M22 S22 G22 S32 S32 NMOS
M32 S32 G32 S42 S42 NMOS
M42 S42 G42 S52 S52 NMOS

M3SSL BL3 G03 S13 S13 NMOS
M13 S13 G13 S23 S23 NMOS
M23 S23 G23 S33 S33 NMOS
M33 S33 G33 S43 S43 NMOS
M43 S43 G43 S53 S53 NMOS

M1SSL BL4 G04 S14 S14 NMOS
M14 S14 G14 S21 S24 NMOS
M24 S24 G24 S34 S34 NMOS
M34 S34 G34 S44 S44 NMOS
M44 S44 G44 S54 S54 NMOS

Look into current comparator.
If current is very small then use current sensing + voltage comparator
