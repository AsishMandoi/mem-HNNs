*NAND_FLASH for Hopfield Network
*A network of 4 transistors in one string and 4 x 5 transistors in x-y plane

Vreadp SL0 gnd 0.5
Vreadn SL1 gnd 0.5
.MODEL NCH0 NMOS LEVEL=72 VERSION=110 BULKMOD=1 GEOMOD=3 L=50n D=10n NBODY=1e21 EOT=28n U0=2e-2 NSD=2e25 RDSMOD=0 PHIG=4.8 RGATEMOD=1 RGEOMOD=1 CGEOMOD=1 RDSW=350 DELVTRAND=677.345m
.MODEL NCH1 NMOS LEVEL=72 VERSION=110 BULKMOD=1 GEOMOD=3 L=50n D=10n NBODY=1e21 EOT=28n U0=2e-2 NSD=2e25 RDSMOD=0 PHIG=4.8 RGATEMOD=1 RGEOMOD=1 CGEOMOD=1 RDSW=350 DELVTRAND=177.345m
.MODEL NCH2 NMOS LEVEL=72 VERSION=110 BULKMOD=1 GEOMOD=3 L=50n D=10n NBODY=1e21 EOT=28n U0=2e-2 NSD=2e25 RDSMOD=0 PHIG=4.8 RGATEMOD=1 RGEOMOD=1 CGEOMOD=1 RDSW=350 DELVTRAND=-322.655m
.MODEL NCH3 NMOS LEVEL=72 VERSION=110 BULKMOD=1 GEOMOD=3 L=50n D=10n NBODY=1e21 EOT=28n U0=2e-2 NSD=2e25 RDSMOD=0 PHIG=4.8 RGATEMOD=1 RGEOMOD=1 CGEOMOD=1 RDSW=350 DELVTRAND=-822.655m
.MODEL NCH4 NMOS LEVEL=72 VERSION=110 BULKMOD=1 GEOMOD=3 L=50n D=10n NBODY=1e21 EOT=28n U0=2e-2 NSD=2e25 RDSMOD=0 PHIG=4.8 RGATEMOD=1 RGEOMOD=1 CGEOMOD=1 RDSW=350 DELVTRAND=-1322.655m
.MODEL NCH5 NMOS LEVEL=72 VERSION=110 BULKMOD=1 GEOMOD=3 L=50n D=10n NBODY=1e21 EOT=28n U0=2e-2 NSD=2e25 RDSMOD=0 PHIG=4.8 RGATEMOD=1 RGEOMOD=1 CGEOMOD=1 RDSW=350 DELVTRAND=-1822.655m
.MODEL NCH6 NMOS LEVEL=72 VERSION=110 BULKMOD=1 GEOMOD=3 L=50n D=10n NBODY=1e21 EOT=28n U0=2e-2 NSD=2e25 RDSMOD=0 PHIG=4.8 RGATEMOD=1 RGEOMOD=1 CGEOMOD=1 RDSW=350 DELVTRAND=-2322.655m
.MODEL NCH7 NMOS LEVEL=72 VERSION=110 BULKMOD=1 GEOMOD=3 L=50n D=10n NBODY=1e21 EOT=28n U0=2e-2 NSD=2e25 RDSMOD=0 PHIG=4.8 RGATEMOD=1 RGEOMOD=1 CGEOMOD=1 RDSW=350 DELVTRAND=-2822.655m
Vselectp G03 gnd 3.5
Vselectn G13 gnd 3.5

VBL01 BL01 gnd 0
VBL11 BL11 gnd 0
VBL02 BL02 gnd 0
VBL12 BL12 gnd 0
VBL03 BL03 gnd 0
VBL13 BL13 gnd 0
VBL04 BL04 gnd 0
VBL14 BL14 gnd 0
VrndPass BSL01 gnd 8
Vpass BSL11 gnd 8
VrndPass BSL02 gnd 0
Vpass BSL12 gnd 8
VrndPass BSL03 gnd 8
Vpass BSL13 gnd 8
VrndPass BSL04 gnd 0
Vpass BSL14 gnd 8
Vpass BSL05 gnd 8
Vpass BSL15 gnd 8



Vpass G02 gnd 8
Vpass G12 gnd 8




Vpass G04 gnd 8
Vpass G14 gnd 8


Vpass G05 gnd 8
Vpass G15 gnd 8



Vpass SSL01 gnd 8
Vpass SSL11 gnd 8
Vpass SSL02 gnd 8
Vpass SSL12 gnd 8
Vpass SSL03 gnd 8
Vpass SSL13 gnd 8
Vpass SSL04 gnd 8
Vpass SSL14 gnd 8
Vpass SSL05 gnd 8
Vpass SSL15 gnd 8

*______+ve Weight Mapping_________

M0111 BL01 BSL01 S0111 S0111 NCH0
M0211 S0111 G02 S0211 S0211 NCH0
M0311 S0211 G03 S0311 S0311 NCH0
M0411 S0311 G04 S0411 S0411 NCH0
M0511 S0411 G05 S0511 S0511 NCH0
M0611 S0511 SSL01 SL0 SL0 NCH0
*One String done
M0121 BL01 BSL02 S0121 S0121 NCH0
M0221 S0121 G02 S0221 S0221 NCH0
M0321 S0221 G03 S0321 S0321 NCH0
M0421 S0321 G04 S0421 S0421 NCH0
M0521 S0421 G05 S0521 S0521 NCH0
M0621 S0521 SSL02 SL0 SL0 NCH0
*One String done
M0131 BL01 BSL03 S0131 S0131 NCH0
M0231 S0131 G02 S0231 S0231 NCH0
M0331 S0231 G03 S0331 S0331 NCH0
M0431 S0331 G04 S0431 S0431 NCH0
M0531 S0431 G05 S0531 S0531 NCH0
M0631 S0531 SSL03 SL0 SL0 NCH0
*One String done
M0141 BL01 BSL04 S0141 S0141 NCH0
M0241 S0141 G02 S0241 S0241 NCH0
M0341 S0241 G03 S0341 S0341 NCH0
M0441 S0341 G04 S0441 S0441 NCH0
M0541 S0441 G05 S0541 S0541 NCH0
M0641 S0541 SSL04 SL0 SL0 NCH0
*One String done
M0151 BL01 BSL05 S0151 S0151 NCH0
M0251 S0151 G02 S0251 S0251 NCH0
M0351 S0251 G03 S0351 S0351 NCH5
M0451 S0351 G04 S0451 S0451 NCH0
M0551 S0451 G05 S0551 S0551 NCH0
M0651 S0551 SSL05 SL0 SL0 NCH0
*One String done
*One yz plane done
M0112 BL02 BSL01 S0112 S0112 NCH0
M0212 S0112 G02 S0212 S0212 NCH0
M0312 S0212 G03 S0312 S0312 NCH0
M0412 S0312 G04 S0412 S0412 NCH0
M0512 S0412 G05 S0512 S0512 NCH0
M0612 S0512 SSL01 SL0 SL0 NCH0
*One String done
M0122 BL02 BSL02 S0122 S0122 NCH0
M0222 S0122 G02 S0222 S0222 NCH0
M0322 S0222 G03 S0322 S0322 NCH0
M0422 S0322 G04 S0422 S0422 NCH0
M0522 S0422 G05 S0522 S0522 NCH0
M0622 S0522 SSL02 SL0 SL0 NCH0
*One String done
M0132 BL02 BSL03 S0132 S0132 NCH0
M0232 S0132 G02 S0232 S0232 NCH0
M0332 S0232 G03 S0332 S0332 NCH0
M0432 S0332 G04 S0432 S0432 NCH0
M0532 S0432 G05 S0532 S0532 NCH0
M0632 S0532 SSL03 SL0 SL0 NCH0
*One String done
M0142 BL02 BSL04 S0142 S0142 NCH0
M0242 S0142 G02 S0242 S0242 NCH0
M0342 S0242 G03 S0342 S0342 NCH0
M0442 S0342 G04 S0442 S0442 NCH0
M0542 S0442 G05 S0542 S0542 NCH0
M0642 S0542 SSL04 SL0 SL0 NCH0
*One String done
M0152 BL02 BSL05 S0152 S0152 NCH0
M0252 S0152 G02 S0252 S0252 NCH0
M0352 S0252 G03 S0352 S0352 NCH5
M0452 S0352 G04 S0452 S0452 NCH0
M0552 S0452 G05 S0552 S0552 NCH0
M0652 S0552 SSL05 SL0 SL0 NCH0
*One String done
*One yz plane done
M0113 BL03 BSL01 S0113 S0113 NCH0
M0213 S0113 G02 S0213 S0213 NCH0
M0313 S0213 G03 S0313 S0313 NCH0
M0413 S0313 G04 S0413 S0413 NCH0
M0513 S0413 G05 S0513 S0513 NCH0
M0613 S0513 SSL01 SL0 SL0 NCH0
*One String done
M0123 BL03 BSL02 S0123 S0123 NCH0
M0223 S0123 G02 S0223 S0223 NCH0
M0323 S0223 G03 S0323 S0323 NCH0
M0423 S0323 G04 S0423 S0423 NCH0
M0523 S0423 G05 S0523 S0523 NCH0
M0623 S0523 SSL02 SL0 SL0 NCH0
*One String done
M0133 BL03 BSL03 S0133 S0133 NCH0
M0233 S0133 G02 S0233 S0233 NCH0
M0333 S0233 G03 S0333 S0333 NCH0
M0433 S0333 G04 S0433 S0433 NCH0
M0533 S0433 G05 S0533 S0533 NCH0
M0633 S0533 SSL03 SL0 SL0 NCH0
*One String done
M0143 BL03 BSL04 S0143 S0143 NCH0
M0243 S0143 G02 S0243 S0243 NCH0
M0343 S0243 G03 S0343 S0343 NCH0
M0443 S0343 G04 S0443 S0443 NCH0
M0543 S0443 G05 S0543 S0543 NCH0
M0643 S0543 SSL04 SL0 SL0 NCH0
*One String done
M0153 BL03 BSL05 S0153 S0153 NCH0
M0253 S0153 G02 S0253 S0253 NCH0
M0353 S0253 G03 S0353 S0353 NCH2
M0453 S0353 G04 S0453 S0453 NCH0
M0553 S0453 G05 S0553 S0553 NCH0
M0653 S0553 SSL05 SL0 SL0 NCH0
*One String done
*One yz plane done
M0114 BL04 BSL01 S0114 S0114 NCH0
M0214 S0114 G02 S0214 S0214 NCH0
M0314 S0214 G03 S0314 S0314 NCH0
M0414 S0314 G04 S0414 S0414 NCH0
M0514 S0414 G05 S0514 S0514 NCH0
M0614 S0514 SSL01 SL0 SL0 NCH0
*One String done
M0124 BL04 BSL02 S0124 S0124 NCH0
M0224 S0124 G02 S0224 S0224 NCH0
M0324 S0224 G03 S0324 S0324 NCH0
M0424 S0324 G04 S0424 S0424 NCH0
M0524 S0424 G05 S0524 S0524 NCH0
M0624 S0524 SSL02 SL0 SL0 NCH0
*One String done
M0134 BL04 BSL03 S0134 S0134 NCH0
M0234 S0134 G02 S0234 S0234 NCH0
M0334 S0234 G03 S0334 S0334 NCH0
M0434 S0334 G04 S0434 S0434 NCH0
M0534 S0434 G05 S0534 S0534 NCH0
M0634 S0534 SSL03 SL0 SL0 NCH0
*One String done
M0144 BL04 BSL04 S0144 S0144 NCH0
M0244 S0144 G02 S0244 S0244 NCH0
M0344 S0244 G03 S0344 S0344 NCH0
M0444 S0344 G04 S0444 S0444 NCH0
M0544 S0444 G05 S0544 S0544 NCH0
M0644 S0544 SSL04 SL0 SL0 NCH0
*One String done
M0154 BL04 BSL05 S0154 S0154 NCH0
M0254 S0154 G02 S0254 S0254 NCH0
M0354 S0254 G03 S0354 S0354 NCH0
M0454 S0354 G04 S0454 S0454 NCH0
M0554 S0454 G05 S0554 S0554 NCH0
M0654 S0554 SSL05 SL0 SL0 NCH0
*One String done
*One yz plane done
*Entire xyz plane done
*______-ve Weight Mapping_________
M1111 BL11 BSL11 S1111 S1111 NCH0
M1211 S1111 G12 S1211 S1211 NCH0
M1311 S1211 G13 S1311 S1311 NCH7
M1411 S1311 G14 S1411 S1411 NCH0
M1511 S1411 G15 S1511 S1511 NCH0
M1611 S1511 SSL11 SL1 SL1 NCH0
*One String done
M1121 BL11 BSL11 S1121 S1121 NCH0
M1221 S1121 G12 S1221 S1221 NCH0
M1321 S1221 G13 S1321 S1321 NCH7
M1421 S1321 G14 S1421 S1421 NCH0
M1521 S1421 G15 S1521 S1521 NCH0
M1621 S1521 SSL12 SL1 SL1 NCH0
*One String done
M1131 BL11 BSL11 S1131 S1131 NCH0
M1231 S1131 G12 S1231 S1231 NCH0
M1331 S1231 G13 S1331 S1331 NCH5
M1431 S1331 G14 S1431 S1431 NCH0
M1531 S1431 G15 S1531 S1531 NCH0
M1631 S1531 SSL13 SL1 SL1 NCH0
*One String done
M1141 BL11 BSL11 S1141 S1141 NCH0
M1241 S1141 G12 S1241 S1241 NCH0
M1341 S1241 G13 S1341 S1341 NCH5
M1441 S1341 G14 S1441 S1441 NCH0
M1541 S1441 G15 S1541 S1541 NCH0
M1641 S1541 SSL14 SL1 SL1 NCH0
*One String done
M1151 BL11 BSL11 S1151 S1151 NCH0
M1251 S1151 G12 S1251 S1251 NCH0
M1351 S1251 G13 S1351 S1351 NCH0
M1451 S1351 G14 S1451 S1451 NCH0
M1551 S1451 G15 S1551 S1551 NCH0
M1651 S1551 SSL15 SL1 SL1 NCH0
*One String done
*One yz plane done
M1112 BL12 BSL11 S1112 S1112 NCH0
M1212 S1112 G12 S1212 S1212 NCH0
M1312 S1212 G13 S1312 S1312 NCH7
M1412 S1312 G14 S1412 S1412 NCH0
M1512 S1412 G15 S1512 S1512 NCH0
M1612 S1512 SSL11 SL1 SL1 NCH0
*One String done
M1122 BL12 BSL11 S1122 S1122 NCH0
M1222 S1122 G12 S1222 S1222 NCH0
M1322 S1222 G13 S1322 S1322 NCH7
M1422 S1322 G14 S1422 S1422 NCH0
M1522 S1422 G15 S1522 S1522 NCH0
M1622 S1522 SSL12 SL1 SL1 NCH0
*One String done
M1132 BL12 BSL11 S1132 S1132 NCH0
M1232 S1132 G12 S1232 S1232 NCH0
M1332 S1232 G13 S1332 S1332 NCH5
M1432 S1332 G14 S1432 S1432 NCH0
M1532 S1432 G15 S1532 S1532 NCH0
M1632 S1532 SSL13 SL1 SL1 NCH0
*One String done
M1142 BL12 BSL11 S1142 S1142 NCH0
M1242 S1142 G12 S1242 S1242 NCH0
M1342 S1242 G13 S1342 S1342 NCH4
M1442 S1342 G14 S1442 S1442 NCH0
M1542 S1442 G15 S1542 S1542 NCH0
M1642 S1542 SSL14 SL1 SL1 NCH0
*One String done
M1152 BL12 BSL11 S1152 S1152 NCH0
M1252 S1152 G12 S1252 S1252 NCH0
M1352 S1252 G13 S1352 S1352 NCH0
M1452 S1352 G14 S1452 S1452 NCH0
M1552 S1452 G15 S1552 S1552 NCH0
M1652 S1552 SSL15 SL1 SL1 NCH0
*One String done
*One yz plane done
M1113 BL13 BSL11 S1113 S1113 NCH0
M1213 S1113 G12 S1213 S1213 NCH0
M1313 S1213 G13 S1313 S1313 NCH5
M1413 S1313 G14 S1413 S1413 NCH0
M1513 S1413 G15 S1513 S1513 NCH0
M1613 S1513 SSL11 SL1 SL1 NCH0
*One String done
M1123 BL13 BSL11 S1123 S1123 NCH0
M1223 S1123 G12 S1223 S1223 NCH0
M1323 S1223 G13 S1323 S1323 NCH5
M1423 S1323 G14 S1423 S1423 NCH0
M1523 S1423 G15 S1523 S1523 NCH0
M1623 S1523 SSL12 SL1 SL1 NCH0
*One String done
M1133 BL13 BSL11 S1133 S1133 NCH0
M1233 S1133 G12 S1233 S1233 NCH0
M1333 S1233 G13 S1333 S1333 NCH7
M1433 S1333 G14 S1433 S1433 NCH0
M1533 S1433 G15 S1533 S1533 NCH0
M1633 S1533 SSL13 SL1 SL1 NCH0
*One String done
M1143 BL13 BSL11 S1143 S1143 NCH0
M1243 S1143 G12 S1243 S1243 NCH0
M1343 S1243 G13 S1343 S1343 NCH0
M1443 S1343 G14 S1443 S1443 NCH0
M1543 S1443 G15 S1543 S1543 NCH0
M1643 S1543 SSL14 SL1 SL1 NCH0
*One String done
M1153 BL13 BSL11 S1153 S1153 NCH0
M1253 S1153 G12 S1253 S1253 NCH0
M1353 S1253 G13 S1353 S1353 NCH0
M1453 S1353 G14 S1453 S1453 NCH0
M1553 S1453 G15 S1553 S1553 NCH0
M1653 S1553 SSL15 SL1 SL1 NCH0
*One String done
*One yz plane done
M1114 BL14 BSL11 S1114 S1114 NCH0
M1214 S1114 G12 S1214 S1214 NCH0
M1314 S1214 G13 S1314 S1314 NCH5
M1414 S1314 G14 S1414 S1414 NCH0
M1514 S1414 G15 S1514 S1514 NCH0
M1614 S1514 SSL11 SL1 SL1 NCH0
*One String done
M1124 BL14 BSL11 S1124 S1124 NCH0
M1224 S1124 G12 S1224 S1224 NCH0
M1324 S1224 G13 S1324 S1324 NCH4
M1424 S1324 G14 S1424 S1424 NCH0
M1524 S1424 G15 S1524 S1524 NCH0
M1624 S1524 SSL12 SL1 SL1 NCH0
*One String done
M1134 BL14 BSL11 S1134 S1134 NCH0
M1234 S1134 G12 S1234 S1234 NCH0
M1334 S1234 G13 S1334 S1334 NCH0
M1434 S1334 G14 S1434 S1434 NCH0
M1534 S1434 G15 S1534 S1534 NCH0
M1634 S1534 SSL13 SL1 SL1 NCH0
*One String done
M1144 BL14 BSL11 S1144 S1144 NCH0
M1244 S1144 G12 S1244 S1244 NCH0
M1344 S1244 G13 S1344 S1344 NCH7
M1444 S1344 G14 S1444 S1444 NCH0
M1544 S1444 G15 S1544 S1544 NCH0
M1644 S1544 SSL14 SL1 SL1 NCH0
*One String done
M1154 BL14 BSL11 S1154 S1154 NCH0
M1254 S1154 G12 S1254 S1254 NCH0
M1354 S1254 G13 S1354 S1354 NCH0
M1454 S1354 G14 S1454 S1454 NCH0
M1554 S1454 G15 S1554 S1554 NCH0
M1654 S1554 SSL15 SL1 SL1 NCH0
*One String done
*One yz plane done
*Entire xyz plane done

OPTION POST=2
PRINT I(VBL01)
PRINT I(VBL02)
.op